// Hello World Test of gowin & the HW-154 Board
