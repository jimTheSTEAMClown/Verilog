// Board configuration: tang_nano_9k_lcd_480_272_tm1638_hackathon
// This module uses few parameterization and relaxed typing rules

module hackathon_top
(
    // System Clocks & Controls  
    input  logic       clock,
    input  logic       slow_clock,
    input  logic       reset,

    // HW-154 I/O Board - Switches & LEDs  
    input  logic [7:0] key,
    output logic [7:0] led,

    // A dynamic seven-segment display  
    output logic [7:0] abcdefgh,
    output logic [7:0] digit,

    // LCD screen interface  
    input  logic [8:0] x,
    input  logic [8:0] y,
    output logic [4:0] red,
    output logic [5:0] green,
    output logic [4:0] blue,

    // HW-154 I/O Board Communication Channel  
    inout  logic [3:0] gpio
);

    //------------------------------------------------------------------------

    // Gates, wires and continuous assignments

    assign led [0] = key [0] & key [1];

    // Exercise 1: Change the code above.
    // Assign to led [0] the result of OR operation (|).

    wire a = key [0];  // Note a new construct - wire
    wire b = key [1];

    assign led [1] = a ^ b; // XOR - eXclusive OR

    //------------------------------------------------------------------------

    
endmodule
